library verilog;
use verilog.vl_types.all;
entity fourBitCounter_vlg_vec_tst is
end fourBitCounter_vlg_vec_tst;
