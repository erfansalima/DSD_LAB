library verilog;
use verilog.vl_types.all;
entity Az1_vlg_check_tst is
    port(
        R3              : in     vl_logic;
        R11             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Az1_vlg_check_tst;
