library verilog;
use verilog.vl_types.all;
entity WaitingRoom_vlg_vec_tst is
end WaitingRoom_vlg_vec_tst;
