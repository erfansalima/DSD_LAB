library verilog;
use verilog.vl_types.all;
entity Az1_vlg_vec_tst is
end Az1_vlg_vec_tst;
